// Code your testbench here
// or browse Examples


module wonscreen(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:29] wonscreen [29:0];
  
  wire [5:0] x = pixel_x[9:4] - 5;
  wire [5:0] y = pixel_y[9:4];
  assign flag = wonscreen[y][x];
  
  initial begin
    wonscreen[0]  = 30'b110110110110110011011011011011; //0
    wonscreen[1]  = 30'b000000000000000000000000000000; //1
    wonscreen[2]  = 30'b000000000000000000000000000000; //2
    wonscreen[3]  = 30'b000000000000000000000000000000; //3
    wonscreen[4]  = 30'b000000000000000000000000000000; //4
    wonscreen[5]  = 30'b010000010000111000010000001000; //5
    wonscreen[6]  = 30'b010000010001000100010000001000; //6
    wonscreen[7]  = 30'b001111100010000010010000001000; //7
    wonscreen[8]  = 30'b000010000100000001010000001000; //8
    wonscreen[9]  = 30'b000010000010000010010000001000; //9
    wonscreen[10] = 30'b000010000001000100010000001000; //10
    wonscreen[11] = 30'b000010000000111000001111110000; //11
    wonscreen[12] = 30'b000000000000000000000000000000; //12
    wonscreen[13] = 30'b000000000000000000000000000000; //13
    wonscreen[14] = 30'b000100000100011100001000000010; //14
    wonscreen[15] = 30'b000100000100100010001100000010; //15
    wonscreen[16] = 30'b000100000101000001001010000010; //16
    wonscreen[17] = 30'b000100000101000001001001000010; //17
    wonscreen[18] = 30'b000100100101000001001000100010; //18
    wonscreen[19] = 30'b000101010101000001001000010010; //19
    wonscreen[20] = 30'b000101010101000001001000001010; //20
    wonscreen[21] = 30'b000110001100100010001000000110; //21
    wonscreen[22] = 30'b000110001100011100001000000010; //22
    wonscreen[23] = 30'b000000000000000000000000000000; //23
    wonscreen[24] = 30'b000000000000000000000000000000; //24
    wonscreen[25] = 30'b000000000000000000000000000000; //25
    wonscreen[26] = 30'b000000000000000000000000000000; //26
    wonscreen[27] = 30'b000000000000000000000000000000; //27
    wonscreen[28] = 30'b000000000000000000000000000000; //28
    wonscreen[29] = 30'b110110110110110011011011011011; //29
  end
endmodule


module startup(pixel_x, pixel_y, squad);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output squad;
  
  reg [0:29] startup [29:0];
  
  wire [5:0] x = pixel_x[9:4] - 5;
  wire [5:0] y = pixel_y[9:4];
  assign squad = startup[y][x];
  
  initial begin
    startup[0]  = 30'b111111111111111111111111111111; 
    startup[1]  = 30'b100000000000000000000000000001; 
    startup[2]  = 30'b100000000000000000000000000001; 
    startup[3]  = 30'b100000000000000000000000000001; 
    startup[4]  = 30'b100000000000000000000000000001; 
    startup[5]  = 30'b100000000000000000000000000001; 
    startup[6]  = 30'b100000000000000000000000000001; 
    startup[7]  = 30'b100000000000000000000000000001; 
    startup[8]  = 30'b100000111011101010111011100001; 
    startup[9]  = 30'b100000100010101010010010100001; 
    startup[10] = 30'b100000111010101010010010100001; 
    startup[11] = 30'b100000001010101010010010100001; 
    startup[12] = 30'b100000001010101010010010100001; 
    startup[13] = 30'b100000111011101110111011100001; 
    startup[14] = 30'b100000000001000000000000000001;
    startup[15] = 30'b100000000000000000000000000001;
    startup[16] = 30'b100000111011101010111011100001; 
    startup[17] = 30'b100000100010101010101010100001; 
    startup[18] = 30'b100000111010101010111010100001; 
    startup[19] = 30'b100000001010101010101010100001; 
    startup[20] = 30'b100000001010101010101010100001; 
    startup[21] = 30'b100000111011101110101011100001; 
    startup[22] = 30'b100000000001000000000000000001; 
    startup[23] = 30'b100000000000000000000000000001; 
    startup[24] = 30'b100000000000000000000000000001; 
    startup[25] = 30'b100000000000000000000000000001; 
    startup[26] = 30'b100000000000000000000000000001; 
    startup[27] = 30'b100000000000000000000000000001; 
    startup[28] = 30'b100000000000000000000000000001; 
    startup[29] = 30'b111111111111111111111111111111; 
  end
endmodule

module lossscreen(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:29] lossscreen [29:0];
  
  wire [5:0] x = pixel_x[9:4] - 5;
  wire [5:0] y = pixel_y[9:4];
  assign flag = lossscreen[y][x];
  
  initial begin
    lossscreen[0]  = 30'b110110110110110011011011011011; //0
    lossscreen[1]  = 30'b000000000000000000000000000000; //1
    lossscreen[2]  = 30'b000000000000000000000000000000; //2
    lossscreen[3]  = 30'b000000000000000000000000000000; //3
    lossscreen[4]  = 30'b000000000000000000000000000000; //4
    lossscreen[5]  = 30'b010000010001110000010000001000; //5
    lossscreen[6]  = 30'b001000100010001000010000001000; //6
    lossscreen[7]  = 30'b000101000100000100010000001000; //7
    lossscreen[8]  = 30'b000010001000000010010000001000; //8
    lossscreen[9]  = 30'b000010000100000100001000001000; //9
    lossscreen[10] = 30'b000010000010001000000100010000; //10
    lossscreen[11] = 30'b000010000001110000000011100000; //11
    lossscreen[12] = 30'b000000000000000000000000000000; //12
    lossscreen[13] = 30'b000000000000000000000000000000; //13
    lossscreen[14] = 30'b010000011110011100001111111100; //14
    lossscreen[15] = 30'b010000010010100000001100000000; //15
    lossscreen[16] = 30'b010000010010100000001100000000; //16
    lossscreen[17] = 30'b010000010010100000001100000000; //17
    lossscreen[18] = 30'b010000010010111100001111110000; //18
    lossscreen[19] = 30'b010000010010000110001100000000; //19
    lossscreen[20] = 30'b010000010010000110001100000000; //20
    lossscreen[21] = 30'b010000010010000110001100000000; //21
    lossscreen[22] = 30'b011111011110111100001111111100; //22
    lossscreen[23] = 30'b000000000000000000000000000000; //23
    lossscreen[24] = 30'b000000000000000000000000000000; //24
    lossscreen[25] = 30'b000000000000000000000000000000; //25
    lossscreen[26] = 30'b000000000000000000000000000000; //26
    lossscreen[27] = 30'b000000000000000000000000000000; //27
    lossscreen[28] = 30'b000000000000000000000000000000; //28
    lossscreen[29] = 30'b110110110110110011011011011011; //29
  end
endmodule



 module red_light(pixel_x, pixel_y, light);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output light;
  
  reg [0:19] red_arr [19:0];
  
   assign light = (((530 <= pixel_x) && (pixel_x< 530 + 20)) && ((110 <= pixel_y) && (pixel_y < 110 + 20))) ? (red_arr[pixel_y - 110][pixel_x - 530]):0;
  initial begin                                      
      red_arr[0]  = 19'b0000000000000000000;   
      red_arr[1]  = 19'b0000000000000000000;   
      red_arr[2]  = 19'b0000000000000000000;    
      red_arr[3]  = 19'b0000000000000000000;   
      red_arr[4]  = 19'b0000011111110000000;   
      red_arr[5]  = 19'b0000111111111100000;   
      red_arr[6]  = 19'b0011111111111110000;   
      red_arr[7]  = 19'b0111111111111111000;   
      red_arr[8]  = 19'b1111111111111111100;   
      red_arr[9]  = 19'b1111111111111111100;   
      red_arr[10] = 19'b1111111111111111100;   
      red_arr[11] = 19'b1111111111111111100;   
      red_arr[12] = 19'b0111111111111111100;   
      red_arr[13] = 19'b0111111111111111000;   
      red_arr[14] = 19'b0011111111111110000;
      red_arr[15] = 19'b0001111111111100000;  
      red_arr[16] = 19'b0000111111110000000;  
      red_arr[17] = 19'b0000000000000000000;  
      red_arr[18] = 19'b0000000000000000000;
      red_arr[19]  = 19'b000000000000000000;      
  end                                                
endmodule
 
 
 module green_light(pixel_x, pixel_y, light);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output light;
  
  reg [0:19] green_arr [19:0];
  
   assign light = (((530 <= pixel_x) && (pixel_x< 530 + 20)) && ((75 <= pixel_y) && (pixel_y < 75 + 20))) ? (green_arr[pixel_y - 75][pixel_x - 530]):0;
  initial begin                                      
      green_arr[0]  = 19'b0000000000000000000;   
      green_arr[1]  = 19'b0000000000000000000;   
      green_arr[2]  = 19'b0000000000000000000;    
      green_arr[3]  = 19'b0000000000000000000;   
      green_arr[4]  = 19'b0000011111110000000;   
      green_arr[5]  = 19'b0000111111111100000;   
      green_arr[6]  = 19'b0011111111111110000;   
      green_arr[7]  = 19'b0111111111111111000;   
      green_arr[8]  = 19'b1111111111111111100;   
      green_arr[9]  = 19'b1111111111111111100;   
      green_arr[10] = 19'b1111111111111111100;   
      green_arr[11] = 19'b1111111111111111100;   
      green_arr[12] = 19'b0111111111111111100;   
      green_arr[13] = 19'b0111111111111111000;   
      green_arr[14] = 19'b0011111111111110000;
      green_arr[15] = 19'b0001111111111100000;  
      green_arr[16] = 19'b0000111111110000000;  
      green_arr[17] = 19'b0000000000000000000;  
      green_arr[18] = 19'b0000000000000000000;
      green_arr[19]  = 19'b000000000000000000;      
  end                                                
endmodule
 
 module maze(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:29] m [29:0];
  
  wire [5:0] x = pixel_x[9:4] - 5;
  wire [5:0] y = pixel_y[9:4];
  assign flag = m[y][x];
  
  initial begin
    m[0]  = 30'b000000000000000000000000000000;
    m[1]  = 30'b111111111100000000001111111111;
    m[2]  = 30'b000000000000000000000000000000;
    m[3]  = 30'b000000000000000000000000111111;
    m[4]  = 30'b000000001000000000000000100000;
    m[5]  = 30'b111111111000000000000000100000;
    m[6]  = 30'b000000000000000000000000000000;
    m[7]  = 30'b000000000000100000000000000000;
    m[8]  = 30'b000000000000111111111110000000;
    m[9]  = 30'b010000001111100000000000000000;
    m[10] = 30'b000000000000100000000000000000;
    m[11] = 30'b111110001111100000000000011111;
    m[12] = 30'b000000000000000000000000000000;
    m[13] = 30'b111111000000000000000000000000;
    m[14] = 30'b000000000000000000100000000000;
    m[15] = 30'b000000000000000000100000000000;
    m[16] = 30'b000000000000011111111000000000;
    m[17] = 30'b000000000000010000000000000000;
    m[18] = 30'b000000000000010000000000000000;
    m[19] = 30'b111100000000010000000000000010;
    m[20] = 30'b000000000000010000000000000010;
    m[21] = 30'b000000000000000000000000000010;
    m[22] = 30'b000000000000000000000000000010;
    m[23] = 30'b011111000000000000000011111110;
    m[24] = 30'b010000000000000000000000000000;
    m[25] = 30'b010000000111111100000000000000;
    m[26] = 30'b010000000000000000000000000000;
    m[27] = 30'b010000000000011110000001110000;
    m[28] = 30'b000000000000000000000000000000;
    m[29] = 30'b000000000000000000000000000000;  
  end
endmodule
 
 module finish(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:19] finish_arr [19:0];
  
   assign flag = (((312 <= pixel_x) && (pixel_x< 312 + 20)) && ((10 <= pixel_y) && (pixel_y < 10 + 20))) ? (finish_arr[pixel_y - 10][pixel_x - 312]):0;
  initial begin                                      
      finish_arr[0]  = 19'b0000000000000000000;   
      finish_arr[1]  = 19'b0000000000000000000;   
      finish_arr[2]  = 19'b1111111111111111100;   
      finish_arr[3]  = 19'b1110000000000000100;  
      finish_arr[4]  = 19'b1110011111111000100;   
      finish_arr[5]  = 19'b1110010000001000100;   
      finish_arr[6]  = 19'b1110010000001000100;   
      finish_arr[7]  = 19'b1110011111111000100;   
      finish_arr[8]  = 19'b1110000000000000100;   
      finish_arr[9]  = 19'b1110000000000000100;   
      finish_arr[10] = 19'b1111111111111111100;   
      finish_arr[11] = 19'b1110000000000000000;   
      finish_arr[12] = 19'b1110000000000000000;   
      finish_arr[13] = 19'b1110000000000000000;   
      finish_arr[14] = 19'b1110000000000000000;   
      finish_arr[15] = 19'b1110000000000000000;
      finish_arr[16] = 19'b1110000000000000000;  
      finish_arr[17] = 19'b0000000000000000000;  
      finish_arr[18] = 19'b0000000000000000000;  
      finish_arr[19] = 19'b0000000000000000000;     
  end                                                
endmodule
 
 module oneheart(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
 reg [0:29] heart_arr [29:0];
  
  
  assign flag = (((450 <= pixel_x) && (pixel_x< 450 + 30)) && ((450 <= pixel_y) && (pixel_y < 450 + 30))) ? (heart_arr[pixel_y - 450][pixel_x - 450]):0;
  
  
  initial begin
    heart_arr[0]  = 30'b000000000000000000000000000000;   
    heart_arr[1]  = 30'b000000000000000000000000000000;   
    heart_arr[2]  = 30'b000000000000000000000000000000;  
    heart_arr[3]  = 30'b000000000000000000000000000000;  
    heart_arr[4]  = 30'b000000000000000000000000000000;    
    heart_arr[5]  = 30'b000000000000000000000000000000;   
    heart_arr[6]  = 30'b000000000000000000000000000000;    
    heart_arr[7]  = 30'b000000000000000000000000000000;    
    heart_arr[8]  = 30'b011101110000000000000000000000;     
    heart_arr[9]  = 30'b111101111000000000000000000000;  
    heart_arr[10] = 30'b011111110000000000000000000000;     
    heart_arr[11] = 30'b001111100000000000000000000000;  
    heart_arr[12] = 30'b000111000000000000000000000000;  
    heart_arr[13] = 30'b000010000000000000000000000000;  
    heart_arr[14] = 30'b000000000000000000000000000000; 
    heart_arr[15] = 30'b000000000000000000000000000000;   
    heart_arr[16] = 30'b000000000000000000000000000000;   
    heart_arr[17] = 30'b000000000000000000000000000000;  
    heart_arr[18] = 30'b000000000000000000000000000000;  
    heart_arr[19] = 30'b000000000000000000000000000000;    
    heart_arr[20] = 30'b000000000000000000000000000000;   
    heart_arr[21] = 30'b000000000000000000000000000000;    
    heart_arr[22] = 30'b000000000000000000000000000000;    
    heart_arr[23] = 30'b000000000000000000000000000000;     
    heart_arr[24] = 30'b000000000000000000000000000000;  
    heart_arr[25] = 30'b000000000000000000000000000000;     
    heart_arr[26] = 30'b000000000000000000000000000000;  
    heart_arr[27] = 30'b000000000000000000000000000000;  
    heart_arr[28] = 30'b000000000000000000000000000000;  
    heart_arr[29] = 30'b000000000000000000000000000000; 
  end
endmodule

module twoheart(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:29] heart_arr [29:0];
  
  
  assign flag = (((450 <= pixel_x) && (pixel_x< 450 + 30)) && ((450 <= pixel_y) && (pixel_y < 450 + 30))) ? (heart_arr[pixel_y - 450][pixel_x - 450]):0;
  
  
  initial begin
    heart_arr[0]  = 30'b000000000000000000000000000000;   
    heart_arr[1]  = 30'b000000000000000000000000000000;   
    heart_arr[2]  = 30'b000000000000000000000000000000;  
    heart_arr[3]  = 30'b000000000000000000000000000000;  
    heart_arr[4]  = 30'b000000000000000000000000000000;    
    heart_arr[5]  = 30'b000000000000000000000000000000;   
    heart_arr[6]  = 30'b000000000000000000000000000000;    
    heart_arr[7]  = 30'b000000000000000000000000000000;    
    heart_arr[8]  = 30'b011101110001110111000000000000;     
    heart_arr[9]  = 30'b111101111011110111100000000000;  
    heart_arr[10] = 30'b011111110001111111000000000000;     
    heart_arr[11] = 30'b001111100000111110000000000000;  
    heart_arr[12] = 30'b000111000000011100000000000000;  
    heart_arr[13] = 30'b000010000000001000000000000000;  
    heart_arr[14] = 30'b000000000000000000000000000000; 
    heart_arr[15] = 30'b000000000000000000000000000000;   
    heart_arr[16] = 30'b000000000000000000000000000000;   
    heart_arr[17] = 30'b000000000000000000000000000000;  
    heart_arr[18] = 30'b000000000000000000000000000000;  
    heart_arr[19] = 30'b000000000000000000000000000000;    
    heart_arr[20] = 30'b000000000000000000000000000000;   
    heart_arr[21] = 30'b000000000000000000000000000000;    
    heart_arr[22] = 30'b000000000000000000000000000000;    
    heart_arr[23] = 30'b000000000000000000000000000000;     
    heart_arr[24] = 30'b000000000000000000000000000000;  
    heart_arr[25] = 30'b000000000000000000000000000000;     
    heart_arr[26] = 30'b000000000000000000000000000000;  
    heart_arr[27] = 30'b000000000000000000000000000000;  
    heart_arr[28] = 30'b000000000000000000000000000000;  
    heart_arr[29] = 30'b000000000000000000000000000000; 
  end
endmodule

module threeheart(pixel_x, pixel_y, flag);
  input [9:0] pixel_x;
  input [9:0] pixel_y;
  output flag;
  
  reg [0:29] heart_arr [29:0];
  
  
  assign flag = (((450 <= pixel_x) && (pixel_x< 450 + 30)) && ((450 <= pixel_y) && (pixel_y < 450 + 30))) ? (heart_arr[pixel_y - 450][pixel_x - 450]):0;

  
  
  initial begin
    heart_arr[0]  = 30'b000000000000000000000000000000;   
    heart_arr[1]  = 30'b000000000000000000000000000000;   
    heart_arr[2]  = 30'b000000000000000000000000000000;  
    heart_arr[3]  = 30'b000000000000000000000000000000;  
    heart_arr[4]  = 30'b000000000000000000000000000000;    
    heart_arr[5]  = 30'b000000000000000000000000000000;   
    heart_arr[6]  = 30'b000000000000000000000000000000;    
    heart_arr[7]  = 30'b000000000000000000000000000000;    
    heart_arr[8]  = 30'b011101110001110111000111011100;     
    heart_arr[9]  = 30'b111101111011110111101111011110;  
    heart_arr[10] = 30'b011111110001111111000111111100;     
    heart_arr[11] = 30'b001111100000111110000011111000;  
    heart_arr[12] = 30'b000111000000011100000001110000;  
    heart_arr[13] = 30'b000010000000001000000000100000;  
    heart_arr[14] = 30'b000000000000000000000000000000; 
    heart_arr[15] = 30'b000000000000000000000000000000;   
    heart_arr[16] = 30'b000000000000000000000000000000;   
    heart_arr[17] = 30'b000000000000000000000000000000;  
    heart_arr[18] = 30'b000000000000000000000000000000;  
    heart_arr[19] = 30'b000000000000000000000000000000;    
    heart_arr[20] = 30'b000000000000000000000000000000;   
    heart_arr[21] = 30'b000000000000000000000000000000;    
    heart_arr[22] = 30'b000000000000000000000000000000;    
    heart_arr[23] = 30'b000000000000000000000000000000;     
    heart_arr[24] = 30'b000000000000000000000000000000;  
    heart_arr[25] = 30'b000000000000000000000000000000;     
    heart_arr[26] = 30'b000000000000000000000000000000;  
    heart_arr[27] = 30'b000000000000000000000000000000;  
    heart_arr[28] = 30'b000000000000000000000000000000;  
    heart_arr[29] = 30'b000000000000000000000000000000; 
  end
endmodule
 
 
module player(clk, ps2_clk, ps2_data, pixel_x, pixel_y, flag, maze_pix, gameend);
  input clk;
  input ps2_clk;
  input ps2_data;
  input [9:0] pixel_x;
  input maze_pix;
  output gameend;
  
  input [9:0] pixel_y;
  reg [3:0]red;
  reg [3:0]green;
  reg [3:0]blue;
  reg [9:0] xpos;
  reg [9:0] ypos;
  reg [3:0] collision = 0;
  reg animate;
  reg gameend;
  reg videoon;

  output flag;
  wire clk_d;
  clk_div_new cd(clk,clk_d);
  wire up, down, left, right, space;
  Keyboard(clk, ps2_clk, ps2_data, up, down, left, right, space);
  
  initial
  begin
  gameend = 0;
  end
  
  
  // initial position of the player
    initial begin
    xpos = 210;
    ypos = 450;
    end
    
    
    //For detecting collission
  
    always @(posedge clk) begin
    if (maze_pix == 1) begin
        if (pixel_y == ypos && ((xpos + 1 <= pixel_x) && (pixel_x<= xpos + 14))) collision[0] = 1;
        if (pixel_y == ypos+15 && ((xpos + 1 <= pixel_x) && (pixel_x< xpos + 14))) collision[1] = 1;
        if (pixel_x == xpos && ((ypos + 1 <= pixel_y) && (pixel_y < ypos + 14))) collision[2] = 1;
        if (pixel_x == xpos+15 && ((ypos + 1 <= pixel_y) && (pixel_y < ypos + 14))) collision[3] = 1;
    
    end
    if (pixel_y == 481 && pixel_x == 0) begin
        collision = 0;
 
    end
    animate <= (pixel_y == 480 && pixel_x == 0); 
  end
  
  // Movement when keys are pressed
  always @(posedge animate) begin
     if (down == 1 && collision[1] == 0) begin
      
        ypos <= ypos + 1;
    
    end
    else if (up == 1 && collision[0] == 0) begin
      
        ypos <= ypos - 1;
     
    end
    else if (left == 1 && collision[2] == 0) begin
        
        xpos <= xpos - 1;
      
    end
    else if (right == 1 && collision[3] == 0) begin
        
        xpos <= xpos + 1;
  
    end
    
    else if(right ==0 && left == 0 && up == 0 && down == 0 && space == 0) begin
    xpos = xpos + 0;
    ypos = ypos + 0;
    end
    
  end
  
  
  //When you reach the finish line, screen switching output goes to pixel gen
  always @(posedge clk)
    begin
    if (ypos <= 30)
    begin
    gameend = 1;
    end
    else
    begin
    gameend = 0;
    end
    end
  
  reg [0:15] m [15:0];
  
   assign flag = (((xpos <= pixel_x) && (pixel_x< xpos + 16)) && ((ypos <= pixel_y) && (pixel_y < ypos + 16))) ? (m[pixel_y - ypos][pixel_x - xpos]):0;
  
  initial begin
    m[0]  = 16'b0000000000000000;
    m[1]  = 16'b0000011111100000;
    m[2]  = 16'b0000111111110000;
    m[3]  = 16'b0001111111111000;
    m[4] =  16'b0011111111111100;
    m[5] =  16'b0011111111111100;
    m[6] =  16'b0111111111111110;
    m[7] =  16'b0100010000100010;
    m[8] =  16'b0100010000100010;
    m[9] =  16'b0110000000000110;
    m[10] = 16'b0010000000000100;
    m[11] = 16'b0011000000001100;
    m[12] = 16'b0001000000001000;
    m[13] = 16'b0001111111111000;
    m[14] = 16'b0000000000000000;
    m[15] = 16'b0000000000000000;  
  end
endmodule
 
 
